module icn (
    input clk_i,
    input rst_i,
    axi_if.Slave  axi_slv,
    axi_if.Master axi_mst
);

endmodule